module  TF_ROM(
    input        [ 7:0] tf_case,
    output logic [22:0] tf_data
);

    always_comb begin
        case(tf_case)
            8'h00:   tf_data = 23'h000001;
            8'h01:   tf_data = 23'h495e02;
            8'h02:   tf_data = 23'h397567;
            8'h03:   tf_data = 23'h396569;
            8'h04:   tf_data = 23'h4f062b;
            8'h05:   tf_data = 23'h53df73;
            8'h06:   tf_data = 23'h4fe033;
            8'h07:   tf_data = 23'h4f066b;
            8'h08:   tf_data = 23'h76b1ae;
            8'h09:   tf_data = 23'h360dd5;
            8'h0a:   tf_data = 23'h28edb0;
            8'h0b:   tf_data = 23'h207fe4;
            8'h0c:   tf_data = 23'h397283;
            8'h0d:   tf_data = 23'h70894a;
            8'h0e:   tf_data = 23'h088192;
            8'h0f:   tf_data = 23'h6d3dc8;
            8'h10:   tf_data = 23'h4c7294;
            8'h11:   tf_data = 23'h41e0b4;
            8'h12:   tf_data = 23'h28a3d2;
            8'h13:   tf_data = 23'h66528a;
            8'h14:   tf_data = 23'h4a18a7;
            8'h15:   tf_data = 23'h794034;
            8'h16:   tf_data = 23'h0a52ee;
            8'h17:   tf_data = 23'h6b7d81;
            8'h18:   tf_data = 23'h4e9f1d;
            8'h19:   tf_data = 23'h1a2877;
            8'h1a:   tf_data = 23'h2571df;
            8'h1b:   tf_data = 23'h1649ee;
            8'h1c:   tf_data = 23'h7611bd;
            8'h1d:   tf_data = 23'h492bb7;
            8'h1e:   tf_data = 23'h2af697;
            8'h1f:   tf_data = 23'h22d8d5;
            8'h20:   tf_data = 23'h36f72a;
            8'h21:   tf_data = 23'h30911e;
            8'h22:   tf_data = 23'h29d13f;
            8'h23:   tf_data = 23'h492673;
            8'h24:   tf_data = 23'h50685f;
            8'h25:   tf_data = 23'h2010a2;
            8'h26:   tf_data = 23'h3887f7;
            8'h27:   tf_data = 23'h11b2c3;
            8'h28:   tf_data = 23'h0603a4;
            8'h29:   tf_data = 23'h0e2bed;
            8'h2a:   tf_data = 23'h10b72c;
            8'h2b:   tf_data = 23'h4a5f35;
            8'h2c:   tf_data = 23'h1f9d15;
            8'h2d:   tf_data = 23'h428cd4;
            8'h2e:   tf_data = 23'h3177f4;
            8'h2f:   tf_data = 23'h20e612;
            8'h30:   tf_data = 23'h341c1d;
            8'h31:   tf_data = 23'h1ad873;
            8'h32:   tf_data = 23'h736681;
            8'h33:   tf_data = 23'h49553f;
            8'h34:   tf_data = 23'h3952f6;
            8'h35:   tf_data = 23'h62564a;
            8'h36:   tf_data = 23'h65ad05;
            8'h37:   tf_data = 23'h439a1c;
            8'h38:   tf_data = 23'h53aa5f;
            8'h39:   tf_data = 23'h30b622;
            8'h3a:   tf_data = 23'h087f38;
            8'h3b:   tf_data = 23'h3b0e6d;
            8'h3c:   tf_data = 23'h2c83da;
            8'h3d:   tf_data = 23'h1c496e;
            8'h3e:   tf_data = 23'h330e2b;
            8'h3f:   tf_data = 23'h1c5b70;
            8'h40:   tf_data = 23'h2ee3f1;
            8'h41:   tf_data = 23'h137eb9;
            8'h42:   tf_data = 23'h57a930;
            8'h43:   tf_data = 23'h3ac6ef;
            8'h44:   tf_data = 23'h3fd54c;
            8'h45:   tf_data = 23'h4eb2ea;
            8'h46:   tf_data = 23'h503ee1;
            8'h47:   tf_data = 23'h7bb175;
            8'h48:   tf_data = 23'h2648b4;
            8'h49:   tf_data = 23'h1ef256;
            8'h4a:   tf_data = 23'h1d90a2;
            8'h4b:   tf_data = 23'h45a6d4;
            8'h4c:   tf_data = 23'h2ae59b;
            8'h4d:   tf_data = 23'h52589c;
            8'h4e:   tf_data = 23'h6ef1f5;
            8'h4f:   tf_data = 23'h3f7288;
            8'h50:   tf_data = 23'h175102;
            8'h51:   tf_data = 23'h075d59;
            8'h52:   tf_data = 23'h1187ba;
            8'h53:   tf_data = 23'h52aca9;
            8'h54:   tf_data = 23'h773e9e;
            8'h55:   tf_data = 23'h0296d8;
            8'h56:   tf_data = 23'h2592ec;
            8'h57:   tf_data = 23'h4cff12;
            8'h58:   tf_data = 23'h404ce8;
            8'h59:   tf_data = 23'h4aa582;
            8'h5a:   tf_data = 23'h1e54e6;
            8'h5b:   tf_data = 23'h4f16c1;
            8'h5c:   tf_data = 23'h1a7e79;
            8'h5d:   tf_data = 23'h03978f;
            8'h5e:   tf_data = 23'h4e4817;
            8'h5f:   tf_data = 23'h31b859;
            8'h60:   tf_data = 23'h5884cc;
            8'h61:   tf_data = 23'h1b4827;
            8'h62:   tf_data = 23'h5b63d0;
            8'h63:   tf_data = 23'h5d787a;
            8'h64:   tf_data = 23'h35225e;
            8'h65:   tf_data = 23'h400c7e;
            8'h66:   tf_data = 23'h6c09d1;
            8'h67:   tf_data = 23'h5bd532;
            8'h68:   tf_data = 23'h6bc4d3;
            8'h69:   tf_data = 23'h258ecb;
            8'h6a:   tf_data = 23'h2e534c;
            8'h6b:   tf_data = 23'h097a6c;
            8'h6c:   tf_data = 23'h3b8820;
            8'h6d:   tf_data = 23'h6d285c;
            8'h6e:   tf_data = 23'h2ca4f8;
            8'h6f:   tf_data = 23'h337caa;
            8'h70:   tf_data = 23'h14b2a0;
            8'h71:   tf_data = 23'h558536;
            8'h72:   tf_data = 23'h28f186;
            8'h73:   tf_data = 23'h55795d;
            8'h74:   tf_data = 23'h4af670;
            8'h75:   tf_data = 23'h234a86;
            8'h76:   tf_data = 23'h75e826;
            8'h77:   tf_data = 23'h78de66;
            8'h78:   tf_data = 23'h05528c;
            8'h79:   tf_data = 23'h7adf59;
            8'h7a:   tf_data = 23'h0f6e17;
            8'h7b:   tf_data = 23'h5bf3da;
            8'h7c:   tf_data = 23'h459b7e;
            8'h7d:   tf_data = 23'h628b34;
            8'h7e:   tf_data = 23'h5dbecb;
            8'h7f:   tf_data = 23'h1a9e7b;
            8'h80:   tf_data = 23'h0006d9;
            8'h81:   tf_data = 23'h6257c5;
            8'h82:   tf_data = 23'h574b3c;
            8'h83:   tf_data = 23'h69a8ef;
            8'h84:   tf_data = 23'h289838;
            8'h85:   tf_data = 23'h64b5fe;
            8'h86:   tf_data = 23'h7ef8f5;
            8'h87:   tf_data = 23'h2a4e78;
            8'h88:   tf_data = 23'h120a23;
            8'h89:   tf_data = 23'h0154a8;
            8'h8a:   tf_data = 23'h09b7ff;
            8'h8b:   tf_data = 23'h435e87;
            8'h8c:   tf_data = 23'h437ff8;
            8'h8d:   tf_data = 23'h5cd5b4;
            8'h8e:   tf_data = 23'h4dc04e;
            8'h8f:   tf_data = 23'h4728af;
            8'h90:   tf_data = 23'h7f735d;
            8'h91:   tf_data = 23'h0c8d0d;
            8'h92:   tf_data = 23'h0f66d5;
            8'h93:   tf_data = 23'h5a6d80;
            8'h94:   tf_data = 23'h61ab98;
            8'h95:   tf_data = 23'h185d96;
            8'h96:   tf_data = 23'h437f31;
            8'h97:   tf_data = 23'h468298;
            8'h98:   tf_data = 23'h662960;
            8'h99:   tf_data = 23'h4bd579;
            8'h9a:   tf_data = 23'h28de06;
            8'h9b:   tf_data = 23'h465d8d;
            8'h9c:   tf_data = 23'h49b0e3;
            8'h9d:   tf_data = 23'h09b434;
            8'h9e:   tf_data = 23'h7c0db3;
            8'h9f:   tf_data = 23'h5a68b0;
            8'ha0:   tf_data = 23'h409ba9;
            8'ha1:   tf_data = 23'h64d3d5;
            8'ha2:   tf_data = 23'h21762a;
            8'ha3:   tf_data = 23'h658591;
            8'ha4:   tf_data = 23'h246e39;
            8'ha5:   tf_data = 23'h48c39b;
            8'ha6:   tf_data = 23'h7bc759;
            8'ha7:   tf_data = 23'h4f5859;
            8'ha8:   tf_data = 23'h392db2;
            8'ha9:   tf_data = 23'h230923;
            8'haa:   tf_data = 23'h12eb67;
            8'hab:   tf_data = 23'h454df2;
            8'hac:   tf_data = 23'h30c31c;
            8'had:   tf_data = 23'h285424;
            8'hae:   tf_data = 23'h13232e;
            8'haf:   tf_data = 23'h7faf80;
            8'hb0:   tf_data = 23'h2dbfcb;
            8'hb1:   tf_data = 23'h022a0b;
            8'hb2:   tf_data = 23'h7e832c;
            8'hb3:   tf_data = 23'h26587a;
            8'hb4:   tf_data = 23'h6b3375;
            8'hb5:   tf_data = 23'h095b76;
            8'hb6:   tf_data = 23'h6be1cc;
            8'hb7:   tf_data = 23'h5e061e;
            8'hb8:   tf_data = 23'h78e00d;
            8'hb9:   tf_data = 23'h628c37;
            8'hba:   tf_data = 23'h3da604;
            8'hbb:   tf_data = 23'h4ae53c;
            8'hbc:   tf_data = 23'h1f1d68;
            8'hbd:   tf_data = 23'h6330bb;
            8'hbe:   tf_data = 23'h7361b8;
            8'hbf:   tf_data = 23'h5ea06c;
            8'hc0:   tf_data = 23'h671ac7;
            8'hc1:   tf_data = 23'h201fc6;
            8'hc2:   tf_data = 23'h5ba4ff;
            8'hc3:   tf_data = 23'h60d772;
            8'hc4:   tf_data = 23'h08f201;
            8'hc5:   tf_data = 23'h6de024;
            8'hc6:   tf_data = 23'h080e6d;
            8'hc7:   tf_data = 23'h56038e;
            8'hc8:   tf_data = 23'h695688;
            8'hc9:   tf_data = 23'h1e6d3e;
            8'hca:   tf_data = 23'h2603bd;
            8'hcb:   tf_data = 23'h6a9dfa;
            8'hcc:   tf_data = 23'h07c017;
            8'hcd:   tf_data = 23'h6dbfd4;
            8'hce:   tf_data = 23'h74d0bd;
            8'hcf:   tf_data = 23'h63e1e3;
            8'hd0:   tf_data = 23'h519573;
            8'hd1:   tf_data = 23'h7ab60d;
            8'hd2:   tf_data = 23'h2867ba;
            8'hd3:   tf_data = 23'h2decd4;
            8'hd4:   tf_data = 23'h58018c;
            8'hd5:   tf_data = 23'h3f4cf5;
            8'hd6:   tf_data = 23'h0b7009;
            8'hd7:   tf_data = 23'h427e23;
            8'hd8:   tf_data = 23'h3cbd37;
            8'hd9:   tf_data = 23'h273333;
            8'hda:   tf_data = 23'h673957;
            8'hdb:   tf_data = 23'h1a4b5d;
            8'hdc:   tf_data = 23'h196926;
            8'hdd:   tf_data = 23'h1ef206;
            8'hde:   tf_data = 23'h11c14e;
            8'hdf:   tf_data = 23'h4c76c8;
            8'he0:   tf_data = 23'h3cf42f;
            8'he1:   tf_data = 23'h7fb19a;
            8'he2:   tf_data = 23'h6af66c;
            8'he3:   tf_data = 23'h2e1669;
            8'he4:   tf_data = 23'h3352d6;
            8'he5:   tf_data = 23'h034760;
            8'he6:   tf_data = 23'h085260;
            8'he7:   tf_data = 23'h741e78;
            8'he8:   tf_data = 23'h2f6316;
            8'he9:   tf_data = 23'h6f0a11;
            8'hea:   tf_data = 23'h07c0f1;
            8'heb:   tf_data = 23'h776d0b;
            8'hec:   tf_data = 23'h0d1ff0;
            8'hed:   tf_data = 23'h345824;
            8'hee:   tf_data = 23'h0223d4;
            8'hef:   tf_data = 23'h68c559;
            8'hf0:   tf_data = 23'h5e8885;
            8'hf1:   tf_data = 23'h2faa32;
            8'hf2:   tf_data = 23'h23fc65;
            8'hf3:   tf_data = 23'h5e6942;
            8'hf4:   tf_data = 23'h51e0ed;
            8'hf5:   tf_data = 23'h65adb3;
            8'hf6:   tf_data = 23'h2ca5e6;
            8'hf7:   tf_data = 23'h79e1fe;
            8'hf8:   tf_data = 23'h7b4064;
            8'hf9:   tf_data = 23'h35e1dd;
            8'hfa:   tf_data = 23'h433aac;
            8'hfb:   tf_data = 23'h464ade;
            8'hfc:   tf_data = 23'h1cfe14;
            8'hfd:   tf_data = 23'h73f1ce;
            8'hfe:   tf_data = 23'h10170e;
            default: tf_data = 23'h74b6d7;
        endcase
    end

endmodule